`timescale 1ns/1ps

//25MHz, %50 duty cycle
module led_blinker #(
    parameter c100 = 125000-1,
    parameter c50  = 250000-1,
    parameter c10  = 1250000-1,
    parameter c1   = 12500000-1
    )(input i_clock, i_enable, i_switch_1, i_switch_2,
    output o_led_drive, dbg_t100, dbg_t50, dbg_t10, dbg_t1, dbg_temp_o_led
);

//en s1 s2 Hz
//0  -  -  -
//1  0  0  100
//1  0  1  50
//1  1  0  10
//1  1  1  1

//keep in mind below that there is 50% duty cycle!
//keep in mind count starts at 0 so do minus 1!
//25MHz = 25,000,000Hz
//100Hz --> count=125,000-1
//50Hz --> count=250,000-1
//10Hz --> count=1,250,000-1
//1Hz --> count=12,500,000-1

//log2(25MHz) --> 25 bits
reg[24:0] count = 0;

//t# = toggle Hz
reg t100 = 1'b0;
reg t50 = 1'b0;
reg t10 = 1'b0;
reg t1 = 1'b0;
reg temp_o_led = 1'b0;

assign dbg_t100 = t100;
assign dbg_t50 = t50;
assign dbg_t10 = t10;
assign dbg_t1 = t1;
assign dbg_temp_o_led = temp_o_led;

// //100hz
// always @(posedge i_clock) begin
     
// end

// //50hz
// always @(posedge i_clock) begin
    
// end

// //10hz
// always @(posedge i_clock) begin
    
// end

// //1hz
// always @(posedge i_clock) begin
    
// end

//count incrementer
always @(posedge i_clock) begin
    if (count>=25000000) begin
        count <= 0;
    end 
    else begin
        count <= count+1;
    end
    if (count%(c100)==0&count!=0) begin
        t100 <= !t100;
    end
    if (count%(c50)==0&count!=0) begin
        t50 <= !t50;
    end 
    if (count%(c10)==0&count!=0) begin
        t10 <= !t10;
    end 
    if (count%(c1)==0&count!=0) begin
        t1 <= !t1;
    end
    if (!i_switch_1&!i_switch_2) begin
        temp_o_led <= t100;
    end else if (!i_switch_1&i_switch_2) begin
        temp_o_led <= t50;
    end else if (i_switch_1&!i_switch_2) begin
        temp_o_led <= t10;
    end else if (i_switch_1&i_switch_2) begin
        temp_o_led <= t1;
    end
end

assign o_led_drive = i_enable & temp_o_led;

endmodule